library verilog;
use verilog.vl_types.all;
entity interface_vlg_vec_tst is
end interface_vlg_vec_tst;
