library verilog;
use verilog.vl_types.all;
entity counter_decoder_vlg_vec_tst is
end counter_decoder_vlg_vec_tst;
