library verilog;
use verilog.vl_types.all;
entity dc_scheme_vlg_vec_tst is
end dc_scheme_vlg_vec_tst;
