library verilog;
use verilog.vl_types.all;
entity scheme1_vlg_vec_tst is
end scheme1_vlg_vec_tst;
