library verilog;
use verilog.vl_types.all;
entity cnteprom_vlg_vec_tst is
end cnteprom_vlg_vec_tst;
