library verilog;
use verilog.vl_types.all;
entity decoder_vlg_check_tst is
    port(
        result          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder_vlg_check_tst;
