library verilog;
use verilog.vl_types.all;
entity counter_logic_vlg_vec_tst is
end counter_logic_vlg_vec_tst;
