library verilog;
use verilog.vl_types.all;
entity speed_loader_vlg_vec_tst is
end speed_loader_vlg_vec_tst;
