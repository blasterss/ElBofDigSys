library verilog;
use verilog.vl_types.all;
entity mux_scheme_vlg_vec_tst is
end mux_scheme_vlg_vec_tst;
