-- megafunction wizard: %LPM_DECODE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_DECODE 

-- ============================================================
-- File Name: lpm_decode3.vhd
-- Megafunction Name(s):
-- 			LPM_DECODE
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.all;

ENTITY lpm_decode3 IS
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
		eq99		: OUT STD_LOGIC 
	);
END lpm_decode3;


ARCHITECTURE SYN OF lpm_decode3 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC ;



	COMPONENT lpm_decode
	GENERIC (
		lpm_decodes		: NATURAL;
		lpm_type		: STRING;
		lpm_width		: NATURAL
	);
	PORT (
			data	: IN STD_LOGIC_VECTOR (6 DOWNTO 0);
			eq	: OUT STD_LOGIC_VECTOR (127 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	sub_wire1    <= sub_wire0(99);
	eq99    <= sub_wire1;

	LPM_DECODE_component : LPM_DECODE
	GENERIC MAP (
		lpm_decodes => 128,
		lpm_type => "LPM_DECODE",
		lpm_width => 7
	)
	PORT MAP (
		data => data,
		eq => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: BaseDec NUMERIC "1"
-- Retrieval info: PRIVATE: EnableInput NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: eq0 NUMERIC "0"
-- Retrieval info: PRIVATE: eq1 NUMERIC "0"
-- Retrieval info: PRIVATE: eq10 NUMERIC "0"
-- Retrieval info: PRIVATE: eq100 NUMERIC "0"
-- Retrieval info: PRIVATE: eq101 NUMERIC "0"
-- Retrieval info: PRIVATE: eq102 NUMERIC "0"
-- Retrieval info: PRIVATE: eq103 NUMERIC "0"
-- Retrieval info: PRIVATE: eq104 NUMERIC "0"
-- Retrieval info: PRIVATE: eq105 NUMERIC "0"
-- Retrieval info: PRIVATE: eq106 NUMERIC "0"
-- Retrieval info: PRIVATE: eq107 NUMERIC "0"
-- Retrieval info: PRIVATE: eq108 NUMERIC "0"
-- Retrieval info: PRIVATE: eq109 NUMERIC "0"
-- Retrieval info: PRIVATE: eq11 NUMERIC "0"
-- Retrieval info: PRIVATE: eq110 NUMERIC "0"
-- Retrieval info: PRIVATE: eq111 NUMERIC "0"
-- Retrieval info: PRIVATE: eq112 NUMERIC "0"
-- Retrieval info: PRIVATE: eq113 NUMERIC "0"
-- Retrieval info: PRIVATE: eq114 NUMERIC "0"
-- Retrieval info: PRIVATE: eq115 NUMERIC "0"
-- Retrieval info: PRIVATE: eq116 NUMERIC "0"
-- Retrieval info: PRIVATE: eq117 NUMERIC "0"
-- Retrieval info: PRIVATE: eq118 NUMERIC "0"
-- Retrieval info: PRIVATE: eq119 NUMERIC "0"
-- Retrieval info: PRIVATE: eq12 NUMERIC "0"
-- Retrieval info: PRIVATE: eq120 NUMERIC "0"
-- Retrieval info: PRIVATE: eq121 NUMERIC "0"
-- Retrieval info: PRIVATE: eq122 NUMERIC "0"
-- Retrieval info: PRIVATE: eq123 NUMERIC "0"
-- Retrieval info: PRIVATE: eq124 NUMERIC "0"
-- Retrieval info: PRIVATE: eq125 NUMERIC "0"
-- Retrieval info: PRIVATE: eq126 NUMERIC "0"
-- Retrieval info: PRIVATE: eq127 NUMERIC "0"
-- Retrieval info: PRIVATE: eq13 NUMERIC "0"
-- Retrieval info: PRIVATE: eq14 NUMERIC "0"
-- Retrieval info: PRIVATE: eq15 NUMERIC "0"
-- Retrieval info: PRIVATE: eq16 NUMERIC "0"
-- Retrieval info: PRIVATE: eq17 NUMERIC "0"
-- Retrieval info: PRIVATE: eq18 NUMERIC "0"
-- Retrieval info: PRIVATE: eq19 NUMERIC "0"
-- Retrieval info: PRIVATE: eq2 NUMERIC "0"
-- Retrieval info: PRIVATE: eq20 NUMERIC "0"
-- Retrieval info: PRIVATE: eq21 NUMERIC "0"
-- Retrieval info: PRIVATE: eq22 NUMERIC "0"
-- Retrieval info: PRIVATE: eq23 NUMERIC "0"
-- Retrieval info: PRIVATE: eq24 NUMERIC "0"
-- Retrieval info: PRIVATE: eq25 NUMERIC "0"
-- Retrieval info: PRIVATE: eq26 NUMERIC "0"
-- Retrieval info: PRIVATE: eq27 NUMERIC "0"
-- Retrieval info: PRIVATE: eq28 NUMERIC "0"
-- Retrieval info: PRIVATE: eq29 NUMERIC "0"
-- Retrieval info: PRIVATE: eq3 NUMERIC "0"
-- Retrieval info: PRIVATE: eq30 NUMERIC "0"
-- Retrieval info: PRIVATE: eq31 NUMERIC "0"
-- Retrieval info: PRIVATE: eq32 NUMERIC "0"
-- Retrieval info: PRIVATE: eq33 NUMERIC "0"
-- Retrieval info: PRIVATE: eq34 NUMERIC "0"
-- Retrieval info: PRIVATE: eq35 NUMERIC "0"
-- Retrieval info: PRIVATE: eq36 NUMERIC "0"
-- Retrieval info: PRIVATE: eq37 NUMERIC "0"
-- Retrieval info: PRIVATE: eq38 NUMERIC "0"
-- Retrieval info: PRIVATE: eq39 NUMERIC "0"
-- Retrieval info: PRIVATE: eq4 NUMERIC "0"
-- Retrieval info: PRIVATE: eq40 NUMERIC "0"
-- Retrieval info: PRIVATE: eq41 NUMERIC "0"
-- Retrieval info: PRIVATE: eq42 NUMERIC "0"
-- Retrieval info: PRIVATE: eq43 NUMERIC "0"
-- Retrieval info: PRIVATE: eq44 NUMERIC "0"
-- Retrieval info: PRIVATE: eq45 NUMERIC "0"
-- Retrieval info: PRIVATE: eq46 NUMERIC "0"
-- Retrieval info: PRIVATE: eq47 NUMERIC "0"
-- Retrieval info: PRIVATE: eq48 NUMERIC "0"
-- Retrieval info: PRIVATE: eq49 NUMERIC "0"
-- Retrieval info: PRIVATE: eq5 NUMERIC "0"
-- Retrieval info: PRIVATE: eq50 NUMERIC "0"
-- Retrieval info: PRIVATE: eq51 NUMERIC "0"
-- Retrieval info: PRIVATE: eq52 NUMERIC "0"
-- Retrieval info: PRIVATE: eq53 NUMERIC "0"
-- Retrieval info: PRIVATE: eq54 NUMERIC "0"
-- Retrieval info: PRIVATE: eq55 NUMERIC "0"
-- Retrieval info: PRIVATE: eq56 NUMERIC "0"
-- Retrieval info: PRIVATE: eq57 NUMERIC "0"
-- Retrieval info: PRIVATE: eq58 NUMERIC "0"
-- Retrieval info: PRIVATE: eq59 NUMERIC "0"
-- Retrieval info: PRIVATE: eq6 NUMERIC "0"
-- Retrieval info: PRIVATE: eq60 NUMERIC "0"
-- Retrieval info: PRIVATE: eq61 NUMERIC "0"
-- Retrieval info: PRIVATE: eq62 NUMERIC "0"
-- Retrieval info: PRIVATE: eq63 NUMERIC "0"
-- Retrieval info: PRIVATE: eq64 NUMERIC "0"
-- Retrieval info: PRIVATE: eq65 NUMERIC "0"
-- Retrieval info: PRIVATE: eq66 NUMERIC "0"
-- Retrieval info: PRIVATE: eq67 NUMERIC "0"
-- Retrieval info: PRIVATE: eq68 NUMERIC "0"
-- Retrieval info: PRIVATE: eq69 NUMERIC "0"
-- Retrieval info: PRIVATE: eq7 NUMERIC "0"
-- Retrieval info: PRIVATE: eq70 NUMERIC "0"
-- Retrieval info: PRIVATE: eq71 NUMERIC "0"
-- Retrieval info: PRIVATE: eq72 NUMERIC "0"
-- Retrieval info: PRIVATE: eq73 NUMERIC "0"
-- Retrieval info: PRIVATE: eq74 NUMERIC "0"
-- Retrieval info: PRIVATE: eq75 NUMERIC "0"
-- Retrieval info: PRIVATE: eq76 NUMERIC "0"
-- Retrieval info: PRIVATE: eq77 NUMERIC "0"
-- Retrieval info: PRIVATE: eq78 NUMERIC "0"
-- Retrieval info: PRIVATE: eq79 NUMERIC "0"
-- Retrieval info: PRIVATE: eq8 NUMERIC "0"
-- Retrieval info: PRIVATE: eq80 NUMERIC "0"
-- Retrieval info: PRIVATE: eq81 NUMERIC "0"
-- Retrieval info: PRIVATE: eq82 NUMERIC "0"
-- Retrieval info: PRIVATE: eq83 NUMERIC "0"
-- Retrieval info: PRIVATE: eq84 NUMERIC "0"
-- Retrieval info: PRIVATE: eq85 NUMERIC "0"
-- Retrieval info: PRIVATE: eq86 NUMERIC "0"
-- Retrieval info: PRIVATE: eq87 NUMERIC "0"
-- Retrieval info: PRIVATE: eq88 NUMERIC "0"
-- Retrieval info: PRIVATE: eq89 NUMERIC "0"
-- Retrieval info: PRIVATE: eq9 NUMERIC "0"
-- Retrieval info: PRIVATE: eq90 NUMERIC "0"
-- Retrieval info: PRIVATE: eq91 NUMERIC "0"
-- Retrieval info: PRIVATE: eq92 NUMERIC "0"
-- Retrieval info: PRIVATE: eq93 NUMERIC "0"
-- Retrieval info: PRIVATE: eq94 NUMERIC "0"
-- Retrieval info: PRIVATE: eq95 NUMERIC "0"
-- Retrieval info: PRIVATE: eq96 NUMERIC "0"
-- Retrieval info: PRIVATE: eq97 NUMERIC "0"
-- Retrieval info: PRIVATE: eq98 NUMERIC "0"
-- Retrieval info: PRIVATE: eq99 NUMERIC "1"
-- Retrieval info: PRIVATE: nBit NUMERIC "7"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_DECODES NUMERIC "128"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DECODE"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "7"
-- Retrieval info: USED_PORT: @eq 0 0 128 0 OUTPUT NODEFVAL "@eq[127..0]"
-- Retrieval info: USED_PORT: data 0 0 7 0 INPUT NODEFVAL "data[6..0]"
-- Retrieval info: USED_PORT: eq99 0 0 0 0 OUTPUT NODEFVAL "eq99"
-- Retrieval info: CONNECT: @data 0 0 7 0 data 0 0 7 0
-- Retrieval info: CONNECT: eq99 0 0 0 0 @eq 0 0 1 99
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode3.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode3.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode3.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode3.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_decode3_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
