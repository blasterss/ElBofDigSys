library verilog;
use verilog.vl_types.all;
entity int_v1_vlg_vec_tst is
end int_v1_vlg_vec_tst;
