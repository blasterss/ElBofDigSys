library verilog;
use verilog.vl_types.all;
entity scheme2_vlg_vec_tst is
end scheme2_vlg_vec_tst;
