library verilog;
use verilog.vl_types.all;
entity count_cycle_vlg_vec_tst is
end count_cycle_vlg_vec_tst;
