library verilog;
use verilog.vl_types.all;
entity prom_mux_vlg_vec_tst is
end prom_mux_vlg_vec_tst;
