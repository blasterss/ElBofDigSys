library verilog;
use verilog.vl_types.all;
entity inter_vlg_vec_tst is
end inter_vlg_vec_tst;
