library verilog;
use verilog.vl_types.all;
entity speed_loader_vlg_check_tst is
    port(
        ModClock        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end speed_loader_vlg_check_tst;
